
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LUT_UN_SIN_128x16 is
	port (
    	phase : in  std_ulogic_vector(6 downto 0);
    	datao : out std_ulogic_vector(15 downto 0) 
  	);
end LUT_UN_SIN_128x16;

architecture lut_arch of LUT_UN_SIN_128x16 is
	type LUT_t is array (natural range 0 to 127) of std_ulogic_vector(15 downto 0);
	constant LUT: LUT_t := (
		0	 =>	 "1000000000000000",
		1	 =>	 "1000011001000111",
		2	 =>	 "1000110010001011",
		3	 =>	 "1001001011000111",
		4	 =>	 "1001100011111000",
		5	 =>	 "1001111100011001",
		6	 =>	 "1010010100100111",
		7	 =>	 "1010101100011111",
		8	 =>	 "1011000011111011",
		9	 =>	 "1011011010111001",
		10	 =>	 "1011110001010110",
		11	 =>	 "1100000111001101",
		12	 =>	 "1100011100011100",
		13	 =>	 "1100110000111111",
		14	 =>	 "1101000100110011",
		15	 =>	 "1101010111110101",
		16	 =>	 "1101101010000010",
		17	 =>	 "1101111011010111",
		18	 =>	 "1110001011110001",
		19	 =>	 "1110011011001111",
		20	 =>	 "1110101001101101",
		21	 =>	 "1110110111001001",
		22	 =>	 "1111000011100010",
		23	 =>	 "1111001110110101",
		24	 =>	 "1111011001000001",
		25	 =>	 "1111100010000100",
		26	 =>	 "1111101001111100",
		27	 =>	 "1111110000101001",
		28	 =>	 "1111110110001001",
		29	 =>	 "1111111010011100",
		30	 =>	 "1111111101100001",
		31	 =>	 "1111111111011000",
		32	 =>	 "1111111111111111",
		33	 =>	 "1111111111011000",
		34	 =>	 "1111111101100001",
		35	 =>	 "1111111010011100",
		36	 =>	 "1111110110001001",
		37	 =>	 "1111110000101001",
		38	 =>	 "1111101001111100",
		39	 =>	 "1111100010000100",
		40	 =>	 "1111011001000001",
		41	 =>	 "1111001110110101",
		42	 =>	 "1111000011100010",
		43	 =>	 "1110110111001001",
		44	 =>	 "1110101001101101",
		45	 =>	 "1110011011001111",
		46	 =>	 "1110001011110001",
		47	 =>	 "1101111011010111",
		48	 =>	 "1101101010000010",
		49	 =>	 "1101010111110101",
		50	 =>	 "1101000100110011",
		51	 =>	 "1100110000111111",
		52	 =>	 "1100011100011100",
		53	 =>	 "1100000111001101",
		54	 =>	 "1011110001010110",
		55	 =>	 "1011011010111001",
		56	 =>	 "1011000011111011",
		57	 =>	 "1010101100011111",
		58	 =>	 "1010010100100111",
		59	 =>	 "1001111100011001",
		60	 =>	 "1001100011111000",
		61	 =>	 "1001001011000111",
		62	 =>	 "1000110010001011",
		63	 =>	 "1000011001000111",
		64	 =>	 "1000000000000000",
		65	 =>	 "0111100110111000",
		66	 =>	 "0111001101110100",
		67	 =>	 "0110110100111000",
		68	 =>	 "0110011100000111",
		69	 =>	 "0110000011100110",
		70	 =>	 "0101101011011000",
		71	 =>	 "0101010011100000",
		72	 =>	 "0100111100000100",
		73	 =>	 "0100100101000110",
		74	 =>	 "0100001110101001",
		75	 =>	 "0011111000110010",
		76	 =>	 "0011100011100011",
		77	 =>	 "0011001111000000",
		78	 =>	 "0010111011001100",
		79	 =>	 "0010101000001010",
		80	 =>	 "0010010101111101",
		81	 =>	 "0010000100101000",
		82	 =>	 "0001110100001110",
		83	 =>	 "0001100100110000",
		84	 =>	 "0001010110010010",
		85	 =>	 "0001001000110110",
		86	 =>	 "0000111100011101",
		87	 =>	 "0000110001001010",
		88	 =>	 "0000100110111110",
		89	 =>	 "0000011101111011",
		90	 =>	 "0000010110000011",
		91	 =>	 "0000001111010110",
		92	 =>	 "0000001001110110",
		93	 =>	 "0000000101100011",
		94	 =>	 "0000000010011110",
		95	 =>	 "0000000000100111",
		96	 =>	 "0000000000000000",
		97	 =>	 "0000000000100111",
		98	 =>	 "0000000010011110",
		99	 =>	 "0000000101100011",
		100	 =>	 "0000001001110110",
		101	 =>	 "0000001111010110",
		102	 =>	 "0000010110000011",
		103	 =>	 "0000011101111011",
		104	 =>	 "0000100110111110",
		105	 =>	 "0000110001001010",
		106	 =>	 "0000111100011101",
		107	 =>	 "0001001000110110",
		108	 =>	 "0001010110010010",
		109	 =>	 "0001100100110000",
		110	 =>	 "0001110100001110",
		111	 =>	 "0010000100101000",
		112	 =>	 "0010010101111101",
		113	 =>	 "0010101000001010",
		114	 =>	 "0010111011001100",
		115	 =>	 "0011001111000000",
		116	 =>	 "0011100011100011",
		117	 =>	 "0011111000110010",
		118	 =>	 "0100001110101001",
		119	 =>	 "0100100101000110",
		120	 =>	 "0100111100000100",
		121	 =>	 "0101010011100000",
		122	 =>	 "0101101011011000",
		123	 =>	 "0110000011100110",
		124	 =>	 "0110011100000111",
		125	 =>	 "0110110100111000",
		126	 =>	 "0111001101110100",
		127	 =>	 "0111100110111000"
  	);
	signal phase_u : unsigned (6 downto 0);

	begin
		phase_u <= unsigned(phase);
		datao <= LUT(to_integer(phase_u)); 
		
end lut_arch;
